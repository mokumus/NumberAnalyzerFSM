module is_odd(
	input  a,
	output o
);

assign o = a;

endmodule